../ccells/s8iom0s8_com_bus_slice_tied_1um.lef